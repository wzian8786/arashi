package arashi_pkg;
    import uvm_pkg::*;

    `include "arashi_param.sv"
    `include "arashi_sequencer.sv"
    `include "arashi_monitor.sv"
    `include "arashi_driver.sv"
    `include "arashi_agent.sv"
    `include "arashi_scoreboard.sv"
    `include "arashi_env.sv"
    `include "arashi_test.sv"
endpackage: arashi_pkg
