`define THREAD_NUM_WIDTH    (2)
`define DATA_WIDTH          (32)
`define MEM_WIDTH           (10)
`define THREAD_NUM          (1 << `THREAD_NUM_WIDTH)
